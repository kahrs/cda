.K DIP2 1 2 -4 -4 4 34
.kp	1 0/0 - 2 0/30

.K DIP8 1 8 -5 0 35 35
.kp	1 0/0 - 4 30/0
.kp	5 30/30 - 8 0/30

.K DIP14 1 14 -9 0 69 31
.kp	1 0/0 - 7 60/0
.kp	8 60/30 - 14 0/30

.K DIP16 1 16 -3 0 73 31
.kp	1 0/0 - 8 70/0
.kp	9 70/30 - 16 0/30

.K LDIP16 1 16 -9 0 79 31
.kp	1 0/0 - 8 70/0
.kp	9 70/30 - 16 0/30

.K DIP18 1 18 -6 0 86 31
.kp	1 0/0 - 9 80/0
.kp	10 80/30 - 18 0/30

.K DIP20 1 20 -6 0 96 31
.kp	1 0/0 - 10 90/0
.kp	11 90/30 - 20 0/30

.K DIP2203 1 22 -5 0 115 31
.kp	1 0/0 - 11 100/0
.kp	12 100/30 - 22 0/30

.K DIP22 1 22 -5 0 115 31
.kp	1 0/0 - 11 100/0
.kp	12 100/30 - 22 0/30

.K DIP2204 1 22 -6 0 106 31
.kp	1 0/0 - 11 100/0
.kp	12 100/40 - 22 0/40

.K DIP2406 1 24 -9 0 119 61
.kp	1 0/0 - 12 110/0
.kp	13 110/60 - 24 0/60

.K DIP24 1 24 -9 0 119 31
.kp	1 0/0 - 12 110/0
.kp	13 110/30 - 24 0/30

.K DIP2403 1 24 -9 0 119 31
.kp	1 0/0 - 12 110/0
.kp	13 110/30 - 24 0/30

.K DIP2404 1 24 -8 0 118 40
.kp	1 0/0 - 12 110/0
.kp	13 110/40 - 24 0/40

.K DIP2806 1 28 -7 0 137 61
.kp	1 0/0 - 14 130/0
.kp	15 130/60 - 28 0/60

.K DIP2804 1 28 -8 -2 138 42
.kp	1 0/0 - 14 130/0
.kp	15 130/40 - 28 0/40

.K DIP2803 1 28 -8 0 138 31
.kp	1 0/0 - 14 130/0
.kp	15 130/30 - 28 0/30

.K DIP28 1 28 -8 0 138 31
.kp	1 0/0 - 14 130/0
.kp	15 130/30 - 28 0/30

.K DIP40 1 40 -9 0 199 61
.kp	1 0/0 - 20 190/0
.kp	21 190/60 - 40 0/60

.K DIP48 1 48 -9 0 239 61
.kp	1 0/0 - 24 230/0
.kp	25 230/60 - 48 0/60

.K DIP48J 1 48 -9 0 239 61
.kp	1 0/0 - 24 230/0
.kp	25 230/60 - 48 0/60

.K DIP64	1 64 -9 0 319 90
.kp	1 0/0 - 32 310/0
.kp	33 310/90 - 64 0/90

.K DIP64J 1 64 -9 0 319 90
.kp	1 0/0 - 32 310/0
.kp	33 310/90 - 64 0/90

.K O4M 1 4 -10 -10 70 40
.kp	1 0/0 - 2 60/0
.kp	3 60/30 - 4 0/30

.K SIP3 1 3 -4 -4 24 4
.kp	1 0/0 - 3 20/0

.K SIP4 1 4 -4 -4 24 4
.kp	1 0/0 - 4 30/0

.K SIP6 1 6 -4 -4 54 4
.kp	1 0/0 - 6 50/0

.K SIP8 1 8 -5 -4 75 4
.kp	1 0/0 - 8 70/0

.K SIP10 1 10 -4 -4 94 4
.kp	1 0/0 - 10 90/0

.K SIP12 1 12 -4 -4 114 4
.kp	1 0/0 - 12 110/0

.K SIP18 1 18 -4 -4 174 4
.kp 1 0/0 - 18 170/0

.K SIP20 1 20 -4 -4 194 4
.kp 1 0/0 - 20 190/0

.K SIP22 1 22 -4 -4 214 4
.kp 1 0/0 - 22 210/0

.K SIP30 1 30 -11 -20 301 -1 %TI mem
.kp	1 0/0 - 30 290/0

.K PG100 1 100 -9 -8 169 108
.kp	1 0/0 - 17 160/0
.kp	18 0/10 - 34 160/10
.kp	35 0/30 - 38 30/30
.kp	39 130/30 - 42 160/30
.kp	43 0/40 - 46 30/40
.kp	47 130/40 - 50 160/40
.kp	51 0/60 - 54 30/60
.kp	55 130/60 - 58 160/60
.kp	59 0/70 - 62 30/70
.kp	63 130/70 - 66 160/70
.kp	67 0/90 - 83 160/90
.kp	84 0/100 - 100 160/100

.K M132 1 132 -9 -8 209 108
.kp	1 0/0 - 21 200/0
.kp	22 0/10 - 42 200/10
.kp	43 0/30 - 48 50/30
.kp	49 150/30 - 54 200/30
.kp	55 0/40 - 60 50/40
.kp	61 150/40 - 66 200/40
.kp	67 0/60 - 72 50/60
.kp	73 150/60 - 78 200/60
.kp	79 0/70 - 84 50/70
.kp	85 150/70 - 90 200/70
.kp	91 0/90 - 111 200/90
.kp	112 0/100 - 132 200/100

.K G114 1 114 -9 -9 129 129	% 68020
.kp 1 0/120 - 13 120/120
.kp 14 0/110 - 26 120/110
.kp 27 0/100 - 39 120/100
.kp 40 0/90 - 42 20/90
.kp 43 110/90 - 44 120/90
.kp 45 0/80 - 47 20/80
.kp 48 110/80 - 49 120/80
.kp 50 0/70 - 52 20/70
.kp 53 110/70 - 54 120/70
.kp 55 0/60 - 57 20/60
.kp 58 100/60 - 60 120/60
.kp 61 0/50 - 63 20/50
.kp 64 110/50 - 65 120/50
.kp 66 0/40 - 68 20/40
.kp 69 110/40 - 70 120/40
.kp 71 0/30 - 73 20/30
.kp 74 110/30 - 75 120/30
.kp 76 0/20 - 88 120/20
.kp 89 0/10 - 101 120/10
.kp 102 0/0 - 114 120/0

.K MG68J 1 68 -9 -9 99 99	% 68881
.kp	1   0/90 - 10 90/90
.kp	11  0/80 - 20 90/80
.kp	21  0/70 - 23 20/70
.kp	24 70/70 - 26 90/70
.kp	27  0/60 - 28 10/60
.kp	29 80/60 - 30 90/60
.kp	31  0/50 - 32 10/50
.kp	33 80/50 - 34 90/50
.kp	35  0/40 - 36 10/40
.kp	37 80/50 - 38 90/40
.kp	39  0/30 - 40 10/30
.kp	41 80/30 - 42 90/30
.kp	43  0/20 - 45 20/20
.kp	46 70/20 - 48 90/20
.kp	49  0/10 - 58 90/10
.kp	59   0/0 - 68 90/0

.K BERG60 1 60 -4 -4 294 14	% Berg
.kd 35
.kp	1 0/0 -2 59 290/0
.kp	2 0/10 -2 60 290/10

.K BERG50 1 50 -4 -4 244 14
.kd 35
.kp	1 0/0 -2 49 240/0
.kp	2 0/10 -2 50 240/10

.K BERG40 1 40 -4 -4 194 14	% Berg
.kd 35
.kp	1 0/0 -2 39 190/0
.kp	2 0/10 -2 40 190/10

.K BERG40R 1 40 -4 -4 196 16 % BERG40 rotated 180
.kd 35
.kp 1 190/0 -2 39 0/0
.kp 2 190/10 -2 40 0/10

.K BERG26 1 26 -4 -4 124 14	% Berg
.kd 35
.kp	1 0/0 -2 25 120/0
.kp	2 0/10 -2 26 120/10

.K BERG20 1 20 -4 -4 94 14	% Berg
.kd 35
.kp	1 0/0 -2 19 90/0
.kp	2 0/10 -2 20 90/10

.K BERG16 1 16 -4 -4 74 14	% Berg
.kd 35
.kp	1 0/0 -2 15 70/0
.kp	2 0/10 -2 16 70/10

.K BERG12 1 12 -4 -4 54 14	% Berg
.kd 35
.kp	1 0/0 -2 11 50/0
.kp	2 0/10 -2 12 50/10

.K BERG10 1 10 -4 -4 44 14	% Berg
.kd 35
.kp	1 0/0 -2 9 40/0
.kp	2 0/10 -2 10 40/10

.K BERG8 1 8 -4 -4 34 14	% Berg
.kd 35
.kp	1 0/0 -2 7 30/0
.kp	2 0/10 -2 8 30/10

.K BERG6 1 6 -4 -4 24 14	% Berg
.kd 35
.kp	1 0/0 -2 5 20/0
.kp	2 0/10 -2 6 20/10

.K DIN96 1 96 -4 -4 24 314
.kd 31
.kp	1 0/0 - 32 0/310
.kp	33 10/0 - 64 10/310
.kp	65 20/0 - 96 20/310

.K PB 1 5 -18 -8 28 28
.kd 40
.kp	1 20/20 - 3 20/0
.kp	4 0/20 - 5 0/0

.K LED 1 2 -4 6 16 -26
.kd 40
.kp	1 0/0 - 2 10/0
